`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NCUT
// Engineer: kayak4665664
// Module Name: prj_30
//////////////////////////////////////////////////////////////////////////////////


module prj_30(
	input [3:0] data,
	output [1:0] out0,
	output [1:0] out1
	);
	assign out0=data[3:2];
	assign out1=data[1:0];
endmodule
