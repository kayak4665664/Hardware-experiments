`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NCUT
// Engineer: kayak4665664
// Module Name: prj_2
//////////////////////////////////////////////////////////////////////////////////

module prj_2(
    input clk,
    output [15:0] sel,
    output [15:0] char
    );
    reg clkout;
    integer cnt;
    integer cnt1;
    reg flag;
    reg [1:0] flag_cnt;
    reg [15:0] scan_cnt;
    parameter period=50;//每一列扫描频率
    parameter sec=15000;//每个字扫描频率
	reg [15:0] ch;
    reg [15:0] s;
    assign char=ch[15:0];//列
    assign sel=s;//片选
    always @(posedge clk)begin//产生扫描频率，控制每一列扫描的快慢
        cnt<=cnt+1;
        if(cnt==(period>>1)-1) clkout<=#1 1'b1;
        else if(cnt==period-1)begin
                clkout<=#1 1'b0;
                cnt<=#1 1'b0;
            end
    end
    always @(posedge clk)begin//产生更换字符的频率，控制每个字扫描的快慢
        cnt1<=cnt1+1;
        if(cnt1==(sec>>1)-1) flag<=#1 1'b1;
        else if(cnt1==sec-1)begin
                flag<=#1 1'b0;
                cnt1<=#1 1'b0;
            end
    end
    always @(posedge clkout)begin//通过扫描频率控制片选和每一列的内容
        scan_cnt<=scan_cnt+1;
        if(scan_cnt=='d15) scan_cnt<=0;
    end
    always @(posedge flag)begin//控制显示的字
        flag_cnt<=flag_cnt+1;
        if(flag_cnt=='d3) flag_cnt<=0;
    end
    always @(scan_cnt)begin
        case(scan_cnt)//片选，选择列
            0:s<=16'b1111111111111110;
            1:s<=16'b1111111111111101;
            2:s<=16'b1111111111111011;
            3:s<=16'b1111111111110111;
            4:s<=16'b1111111111101111;
            5:s<=16'b1111111111011111;
            6:s<=16'b1111111110111111;
            7:s<=16'b1111111101111111;
            8:s<=16'b1111111011111111;
            9:s<=16'b1111110111111111;
            10:s<=16'b1111101111111111;
            11:s<=16'b1111011111111111;
            12:s<=16'b1110111111111111;
            13:s<=16'b1101111111111111;
            14:s<=16'b1011111111111111;
            15:s<=16'b0111111111111111;
            default:s<=16'b1111111111111111;
        endcase
    end
    always @(scan_cnt)begin
        if(!flag_cnt)
            case(scan_cnt)//X
                0:ch=16'b0000000000000000;
                1:ch=16'b0000000000000000;
                2:ch=16'b0000000000000000;
                3:ch=16'b0000000000000000;
                4:ch=16'b0000000000000000;
                5:ch=16'b0000000000000000;
                6:ch=16'b0000000000000000;
                7:ch=16'b0000000000000000;
                8:ch=16'b0000000000000000;
                9:ch=16'b0000000000000000;
                10:ch=16'b0000000000000000;
                11:ch=16'b0000000000000000;
                12:ch=16'b0000000000000000;
                13:ch=16'b0000000000000000;
                14:ch=16'b0000000000000000;
                15:ch=16'b0000000000000000;
                default:ch=16'b0000000000000000;
            endcase
        else if(flag_cnt==1||flag_cnt==3)
            case(scan_cnt)//X
                0:ch=16'b0000000000000000;
                1:ch=16'b0000000000000000;
                2:ch=16'b0000000000000000;
                3:ch=16'b0000000000000000;
                4:ch=16'b0000000000000000;
                5:ch=16'b0000000000000000;
                6:ch=16'b0000000000000000;
                7:ch=16'b0000000000000000;
                8:ch=16'b0000000000000000;
                9:ch=16'b0000000000000000;
                10:ch=16'b0000000000000000;
                11:ch=16'b0000000000000000;
                12:ch=16'b0000000000000000;
                13:ch=16'b0000000000000000;
                14:ch=16'b0000000000000000;
                15:ch=16'b0000000000000000;
                default:ch=16'b0000000000000000;
            endcase
        else
            case(scan_cnt)//X
                0:ch=16'b0000000000000000;
                1:ch=16'b0000000000000000;
                2:ch=16'b0000000000000000;
                3:ch=16'b0000000000000000;
                4:ch=16'b0000000000000000;
                5:ch=16'b0000000000000000;
                6:ch=16'b0000000000000000;
                7:ch=16'b0000000000000000;
                8:ch=16'b0000000000000000;
                9:ch=16'b0000000000000000;
                10:ch=16'b0000000000000000;
                11:ch=16'b0000000000000000;
                12:ch=16'b0000000000000000;
                13:ch=16'b0000000000000000;
                14:ch=16'b0000000000000000;
                15:ch=16'b0000000000000000;
                default:ch=16'b0000000000000000;
            endcase
    end
endmodule